library verilog;
use verilog.vl_types.all;
entity mips_single_cycle_tb is
end mips_single_cycle_tb;
