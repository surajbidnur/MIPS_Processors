library verilog;
use verilog.vl_types.all;
entity mips_multi_cycle_tb is
end mips_multi_cycle_tb;
