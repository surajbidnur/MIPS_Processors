library verilog;
use verilog.vl_types.all;
entity mips_pipeline_processor_tb is
end mips_pipeline_processor_tb;
